module absdb(
  input [0:127] ra,
  input [0:127] rb,

  output reg [0:127] result
);
integer j;

always @(*) begin
  for (j = 0; j < 16; j = j + 1) begin
    if (ra[8*j +: 8] < rb[8*j +: 8]) begin
      result[8*j +: 8] = rb[8*j +: 8] - ra[8*j +: 8];
    end else begin
      result[8*j +: 8] = ra[8*j +: 8] - rb[8*j +: 8];
    end
  end
end

endmodule