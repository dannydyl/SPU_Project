module Decode_HzdCheck(
  input clk,
  input rst,
  input [0:31] instruction_in1,
  input [0:31] instruction_in2,


);

endmodule