module Decode_HzdCheck(
  input clk,
  input rst,
  input [31:0] instruction_in1,
  input [31:0] instruction_in2,

  
);

endmodule